
program main();


   import uvm_pkg::*;

   `include "testcase1.sv"

   initial begin
   
      run_test(); // uvm_top.run_test();

   end

endprogram


